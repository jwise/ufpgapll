module IBUFG(output wire O, input I);
  assign O = I;
endmodule
